module adder(r,s,u);
input [31:0] r,s;
output [31:0] u;
assign u = r+s;
endmodule
